`ifndef MEMORY_PKG_SV
 `define MEMORY_PKG_SV

package memory_pkg;

 `include "v2_tr.sv"
 `include "v2_driver.sv"
 `include "v2_monitor.sv"

endpackage : memory_pkg

`endif
